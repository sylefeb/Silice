`define FORMAL 1
$$NUM_LEDS=8

module top();
// do nothing
endmodule
