module differential_pair(
        input  I,
        output OT,
        output OC
    );

OBCO dp(.I(I), .OT(OT), .OC(OC) );

endmodule
