module vfoo(input [7:0] v,output [7:0] o);

  assign o = v;

endmodule
